/************************************************************
* Filename      : chiplet.sv
* Author        : kiki
* Create        : 2023-03-10 09:23:40
* Last Modified : 2023-03-14 09:08:49
* Description   : This is a production script.
************************************************************/

module chiplet(
input               pad18_xin_osc,
input               pad18_po_reset_n,
input       [1:0]   pad18_chip_mode,
input       [2:0]   pad18_my_chip_x,
input       [2:0]   pad18_my_chip_y,
input       [7:0]   pad18_cfg_io,
inout  wire [31:0]  pad18_gpio,
input               pad18_uart0_rx_i,
output wire         pad18_uart0_tx_o,
input               pad18_uart1_rx_i,
output wire         pad18_uart1_tx_o,
input               pad18_spi_s0_clk_i,
input               pad18_spi_s0_cs_i,
output wire         pad18_spi_s0_sdo0_o,
input               pad18_spi_s0_sdi0_i,
input               pad18_spi_s1_clk_i,
input               pad18_spi_s1_cs_i,
output wire         pad18_spi_s1_sdo0_o,
input               pad18_spi_s1_sdi0_i,
output wire         pad18_spi_m_clk_o,
output wire         pad18_spi_m_csn0_o,
output wire         pad18_spi_m_csn1_o,
output wire         pad18_spi_m_csn2_o,
output wire         pad18_spi_m_csn3_o,
output wire         pad18_spi_m_sdo0_o,
input               pad18_spi_m_sdi0_i,
inout  wire         pad18_scl,
inout  wire         pad18_sda,
input               pad18_tck_i,
input               pad18_trstn_i,
input               pad18_tms_i,
input               pad18_tdi_i,
output wire         pad18_tdo_o,
inout  wire [31:0]  pad18_sdram_data,
output wire [3:0]   pad18_sdram_dqm,
output wire [3:0]   pad18_sdram_cs_n_o,
output wire [14:0]  pad18_sdram_addr_o,
output wire [3:0]   pad18_sdram_cke_o,
output wire         pad18_sdram_ras_n_o,
output wire         pad18_sdram_cas_n_o,
output wire         pad18_sdram_we_n_o,
output wire         pad18_sdram_clk_o,
output wire         pada_pll_atest0,
output wire         pada_pll_atest1,
input       [9:0]   pad18_dbg_mux_cfg,
output wire         pad18_test_signal_out,
output wire         pad09_east_dcc_atb,
output wire         pad09_west_dcc_atb,
output wire         pad09_north_dcc_atb,
output wire         pad09_south_dcc_atb,
output wire [79:0]  pad09_east_tx,
input       [79:0]  pad09_east_rx,
output wire         pad09_east_ns_fwd_clk,
output wire         pad09_east_ns_fwd_clkb,
output wire         pad09_east_ns_sr_clk,
output wire         pad09_east_ns_sr_clkb,
output wire         pad09_east_ns_sr_load,
output wire         pad09_east_ns_sr_data,
output wire         pad09_east_ns_mac_rdy,
output wire         pad09_east_ns_adapter_rstn,
output wire         pad09_east_spare1_out,
output wire         pad09_east_spare0_out,
input               pad09_east_fs_fwd_clk,
input               pad09_east_fs_fwd_clkb,
input               pad09_east_fs_sr_clk,
input               pad09_east_fs_sr_clkb,
input               pad09_east_fs_sr_load,
input               pad09_east_fs_sr_data,
input               pad09_east_fs_mac_rdy,
input               pad09_east_fs_adapter_rstn,
input               pad09_east_spare1_in,
input               pad09_east_spare0_in,
output wire [79:0]  pad09_south_tx,
input       [79:0]  pad09_south_rx,
output wire         pad09_south_ns_fwd_clk,
output wire         pad09_south_ns_fwd_clkb,
output wire         pad09_south_ns_sr_clk,
output wire         pad09_south_ns_sr_clkb,
output wire         pad09_south_ns_sr_load,
output wire         pad09_south_ns_sr_data,
output wire         pad09_south_ns_mac_rdy,
output wire         pad09_south_ns_adapter_rstn,
output wire         pad09_south_spare1_out,
output wire         pad09_south_spare0_out,
input               pad09_south_fs_fwd_clkb,
input               pad09_south_fs_fwd_clk,
input               pad09_south_fs_sr_clkb,
input               pad09_south_fs_sr_clk,
input               pad09_south_fs_sr_load,
input               pad09_south_fs_sr_data,
input               pad09_south_fs_mac_rdy,
input               pad09_south_fs_adapter_rstn,
input               pad09_south_spare1_in,
input               pad09_south_spare0_in,
output wire [79:0]  pad09_west_tx,
input       [79:0]  pad09_west_rx,
output wire         pad09_west_ns_fwd_clk,
output wire         pad09_west_ns_fwd_clkb,
output wire         pad09_west_ns_sr_clk,
output wire         pad09_west_ns_sr_clkb,
output wire         pad09_west_ns_sr_load,
output wire         pad09_west_ns_sr_data,
output wire         pad09_west_ns_mac_rdy,
output wire         pad09_west_ns_adapter_rstn,
output wire         pad09_west_spare1_out,
output wire         pad09_west_spare0_out,
input               pad09_west_fs_fwd_clkb,
input               pad09_west_fs_fwd_clk,
input               pad09_west_fs_sr_clkb,
input               pad09_west_fs_sr_clk,
input               pad09_west_fs_sr_load,
input               pad09_west_fs_sr_data,
input               pad09_west_fs_mac_rdy,
input               pad09_west_fs_adapter_rstn,
input               pad09_west_spare1_in,
input               pad09_west_spare0_in,
output wire [79:0]  pad09_north_tx,
input       [79:0]  pad09_north_rx,
output wire         pad09_north_ns_fwd_clk,
output wire         pad09_north_ns_fwd_clkb,
output wire         pad09_north_ns_sr_clk,
output wire         pad09_north_ns_sr_clkb,
output wire         pad09_north_ns_sr_load,
output wire         pad09_north_ns_sr_data,
output wire         pad09_north_ns_mac_rdy,
output wire         pad09_north_ns_adapter_rstn,
output wire         pad09_north_spare1_out,
output wire         pad09_north_spare0_out,
input               pad09_north_fs_fwd_clkb,
input               pad09_north_fs_fwd_clk,
input               pad09_north_fs_sr_clkb,
input               pad09_north_fs_sr_clk,
input               pad09_north_fs_sr_load,
input               pad09_north_fs_sr_data,
input               pad09_north_fs_mac_rdy,
input               pad09_north_fs_adapter_rstn,
input               pad09_north_spare1_in,
input               pad09_north_spare0_in
);


endmodule


`endif
